LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.all;
PACKAGE data_maps IS
type maps_type is array (1 to 22,1 to 23) of integer range 0 to 5;
END data_maps;