LIBRARY IEEE;
USE  IEEE.STD_LOGIC_1164.all;
USE IEEE.STD_LOGIC_ARITH.all;
USE  IEEE.STD_LOGIC_UNSIGNED.all;

ENTITY Char_ROM IS
	PORT(	character_address		: 	IN	STD_LOGIC_VECTOR(7 DOWNTO 0);
			font_row, font_col		: 	IN 	STD_LOGIC_VECTOR(2 DOWNTO 0);
			rom_mux_output			: 	OUT	STD_LOGIC);
END Char_ROM;

ARCHITECTURE a OF Char_ROM IS
	SIGNAL	rom_data			: STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL	rom_address			: STD_LOGIC_VECTOR(10 DOWNTO 0);
BEGIN
				-- Small 8 by 8 Character Generator ROM for Video Display
				-- Each character is eight 8-bits words of pixel data
With rom_address select
				--@
	rom_data <= "00111100" 	when "01000000000",
				"01100110" 	when "01000000001",
				"01101110" 	when "01000000010",
				"01101110" 	when "01000000011",
				"01100000" 	when "01000000100",
				"01100010" 	when "01000000101",
	 			"00111100" 	when "01000000110",
				"00000000" 	when "01000000111",
				--A
				"00011000"	when "01000001000",
				"00111100"	when "01000001001",
				"01100110"	when "01000001010",
				"01111110"	when "01000001011",
				"01100110"	when "01000001100",
				"01100110"	when "01000001101",
				"01100110"	when "01000001110",
				"00000000"	when "01000001111",
				--B
				"01111100" 	when "01000010000",
				"01100110" 	when "01000010001",
				"01100110" 	when "01000010010",
				"01111100" 	when "01000010011",
				"01100110" 	when "01000010100",
				"01100110" 	when "01000010101",
	 			"01111100" 	when "01000010110",
				"00000000"	when "01000010111",				

				--C
				"00111100" 	when "01000011000",
				"01100110" 	when "01000011001",
				"01100000" 	when "01000011010",
				"01100000" 	when "01000011011",
				"01100000" 	when "01000011100",
				"01100110" 	when "01000011101",
	 			"00111100" 	when "01000011110",
				"00000000"	when "01000011111",
				--D
				"01111000" 	when "01000100000",
				"01101100" 	when "01000100001",
				"01100110" 	when "01000100010",
				"01100110" 	when "01000100011",
				"01100110" 	when "01000100100",
				"01101100" 	when "01000100101",
	 			"01111000" 	when "01000100110",
				"00000000"	when "01000100111",				

				--E
				"01111110" 	when "01000101000",
				"01100000" 	when "01000101001",
				"01100000" 	when "01000101010",
				"01111000" 	when "01000101011",
				"01100000" 	when "01000101100",
				"01100000" 	when "01000101101",
	 			"01111110" 	when "01000101110",
				"00000000"	when "01000101111",
				--F
				"01111110" 	when "01000110000",--0
				"01100000" 	when "01000110001",--1
				"01100000" 	when "01000110010",--2
				"01111000" 	when "01000110011",--3
				"01100000" 	when "01000110100",--4
				"01100000" 	when "01000110101",--5
	 			"01100000" 	when "01000110110",--6
				"00000000"	when "01000110111",--7
				--G
				"00111100" 	when "01000111000",--0
				"01100110" 	when "01000111001",--1
				"01100000" 	when "01000111010",--2
				"01101110" 	when "01000111011",--3
				"01100110" 	when "01000111100",--4
				"01100110" 	when "01000111101",--5
	 			"00111100" 	when "01000111110",--6
				"00000000"	when "01000111111",--7
				--H
				"01100110" 	when "01001000000",--0
				"01100110" 	when "01001000001",--1
				"01100110" 	when "01001000010",--2
				"01111110" 	when "01001000011",--3
				"01100110" 	when "01001000100",--4
				"01100110" 	when "01001000101",--5
	 			"01100110" 	when "01001000110",--6
				"00000000"	when "01001000111",--7
				--I
				"00111100" 	when "01001001000",--0
				"00011000" 	when "01001001001",--1
				"00011000" 	when "01001001010",--2
				"00011000" 	when "01001001011",--3
				"00011000" 	when "01001001100",--4
				"00011000" 	when "01001001101",--5
	 			"00111100" 	when "01001001110",--6
				"00000000"	when "01001001111",--7
				--J
				"00011110" 	when "01001010000",--0
				"00001100" 	when "01001010001",--1
				"00001100" 	when "01001010010",--2
				"00001100" 	when "01001010011",--3
				"00001100" 	when "01001010100",--4
				"01101100" 	when "01001010101",--5
	 			"00111000" 	when "01001010110",--6
				"00000000"	when "01001010111",--7
				--K
				"01100110" 	when "01001011000",--0
				"01101100" 	when "01001011001",--1
				"01111000" 	when "01001011010",--2
				"01110000" 	when "01001011011",--3
				"01111000" 	when "01001011100",--4
				"01101100" 	when "01001011101",--5
	 			"01100110" 	when "01001011110",--6
				"00000000"	when "01001011111",--7
				--L
				"01100000" 	when "01001100000",--0
				"01100000" 	when "01001100001",--1
				"01100000" 	when "01001100010",--2
				"01100000" 	when "01001100011",--3
				"01100000" 	when "01001100100",--4
				"01100000" 	when "01001100101",--5
	 			"01111110" 	when "01001100110",--6
				"00000000"	when "01001100111",--7
				--M
				"01100011" 	when "01001101000",--0
				"01110111" 	when "01001101001",--1
				"01111111" 	when "01001101010",--2
				"01101011" 	when "01001101011",--3
				"01100011" 	when "01001101100",--4
				"01100011" 	when "01001101101",--5
	 			"01100011" 	when "01001101110",--6
				"00000000"	when "01001101111",--7
				--N
				"01100110" 	when "01001110000",--0
				"01100110" 	when "01001110001",--1
				"01111110" 	when "01001110010",--2
				"01111110" 	when "01001110011",--3
				"01101110" 	when "01001110100",--4
				"01100110" 	when "01001110101",--5
	 			"01100110" 	when "01001110110",--6
				"00000000"	when "01001110111",--7
				--O
				"00111100" 	when "01001111000",--0
				"01100110" 	when "01001111001",--1
				"01100110" 	when "01001111010",--2
				"01100110" 	when "01001111011",--3
				"01100110" 	when "01001111100",--4
				"01100110" 	when "01001111101",--5
	 			"00111100" 	when "01001111110",--6
				"00000000"	when "01001111111",--7
				--P
				"01111100" 	when "01010000000",--0
				"01100110" 	when "01010000001",--1
				"01100110" 	when "01010000010",--2
				"01111100" 	when "01010000011",--3
				"01100000" 	when "01010000100",--4
				"01100000" 	when "01010000101",--5
	 			"01100000" 	when "01010000110",--6
				"00000000"	when "01010000111",--7
				--Q
				"00111100" 	when "01010001000",--0
				"01100110" 	when "01010001001",--1
				"01100110" 	when "01010001010",--2
				"01100110" 	when "01010001011",--3
				"01100110" 	when "01010001100",--4
				"00111100" 	when "01010001101",--5
	 			"00001110" 	when "01010001110",--6
				"00000000"	when "01010001111",--7
				--R
				"01111100" 	when "01010010000",--0
				"01100110" 	when "01010010001",--1
				"01100110" 	when "01010010010",--2
				"01111100" 	when "01010010011",--3
				"01111000" 	when "01010010100",--4
				"01101100" 	when "01010010101",--5
	 			"01100110" 	when "01010010110",--6
				"00000000"	when "01010010111",--7
				--S
				"00111100" 	when "01010011000",--0
				"01100110" 	when "01010011001",--1
				"01100000" 	when "01010011010",--2
				"00111100" 	when "01010011011",--3
				"00000110" 	when "01010011100",--4
				"01100110" 	when "01010011101",--5
	 			"00111100" 	when "01010011110",--6
				"00000000"	when "01010011111",--7
				--T
				"01111110" 	when "01010100000",--0
				"00011000" 	when "01010100001",--1
				"00011000" 	when "01010100010",--2
				"00011000" 	when "01010100011",--3
				"00011000" 	when "01010100100",--4
				"00011000" 	when "01010100101",--5
	 			"00011000" 	when "01010100110",--6
				"00000000"	when "01010100111",--7
				--U
				"01100110" 	when "01010101000",--0
				"01100110" 	when "01010101001",--1
				"01100110" 	when "01010101010",--2
				"01100110" 	when "01010101011",--3
				"01100110" 	when "01010101100",--4
				"01100110" 	when "01010101101",--5
	 			"00111100" 	when "01010101110",--6
				"00000000"	when "01010101111",--7
				--V
				"01100110" 	when "01010110000",--0
				"01100110" 	when "01010110001",--1
				"01100110" 	when "01010110010",--2
				"01100110" 	when "01010110011",--3
				"01100110" 	when "01010110100",--4
				"00111100" 	when "01010110101",--5
	 			"00011000" 	when "01010110110",--6
				"00000000"	when "01010110111",--7
				--W
				"01100011" 	when "01010111000",--0
				"01100011" 	when "01010111001",--1
				"01100011" 	when "01010111010",--2
				"01101011" 	when "01010111011",--3
				"01111111" 	when "01010111100",--4
				"01110111" 	when "01010111101",--5
	 			"01100011" 	when "01010111110",--6
				"00000000"	when "01010111111",--7
				--X
				"01100110" 	when "01011000000",--0
				"01100110" 	when "01011000001",--1
				"00111100" 	when "01011000010",--2
				"00011000" 	when "01011000011",--3
				"00111100" 	when "01011000100",--4
				"01100110" 	when "01011000101",--5
	 			"01100110" 	when "01011000110",--6
				"00000000"	when "01011000111",--7
				--Y
				"01100110" 	when "01011001000",--0
				"01100110" 	when "01011001001",--1
				"01100110" 	when "01011001010",--2
				"00111100" 	when "01011001011",--3
				"00011000" 	when "01011001100",--4
				"00011000" 	when "01011001101",--5
	 			"00011000" 	when "01011001110",--6
				"00000000"	when "01011001111",--7
				--Z
				"01111110" 	when "01011010000",--0
				"00000110" 	when "01011010001",--1
				"00001100" 	when "01011010010",--2
				"00011000" 	when "01011010011",--3
				"00110000" 	when "01011010100",--4
				"01100000" 	when "01011010101",--5
	 			"01111110" 	when "01011010110",--6
				"00000000"	when "01011010111",--7
				--[
				"00111100" 	when "01011011000",--0
				"00110000" 	when "01011011001",--1
				"00110000" 	when "01011011010",--2
				"00110000" 	when "01011011011",--3
				"00110000" 	when "01011011100",--4
				"00110000" 	when "01011011101",--5
	 			"00111100" 	when "01011011110",--6
				"00000000"	when "01011011111",--7
				--\--
				"00000000" 	when "01011100000",--0
				"11000000" 	when "01011100001",--1
				"01100000" 	when "01011100010",--2
				"00110000" 	when "01011100011",--3
				"00011000" 	when "01011100100",--4
				"00001100" 	when "01011100101",--5
	 			"00000110" 	when "01011100110",--6
				"00000000"	when "01011100111",--7
				--]
				"00111100" 	when "01011101000",--0
				"00001100" 	when "01011101001",--1
				"00001100" 	when "01011101010",--2
				"00001100" 	when "01011101011",--3
				"00001100" 	when "01011101100",--4
				"00001100" 	when "01011101101",--5
	 			"00111100" 	when "01011101110",--6
				"00000000"	when "01011101111",--7
				--^
				"00000000" 	when "01011110000",--0
				"00011000" 	when "01011110001",--1
				"00111100" 	when "01011110010",--2
				"01100110" 	when "01011110011",--3
				"00000000" 	when "01011110100",--4
				"00000000" 	when "01011110101",--5
	 			"00000000" 	when "01011110110",--6
				"00000000"	when "01011110111",--7
				--_
				"00000000" 	when "01011111000",--0
				"00000000" 	when "01011111001",--1
				"00000000" 	when "01011111010",--2
				"00000000" 	when "01011111011",--3
				"00000000" 	when "01011111100",--4
				"00000000" 	when "01011111101",--5
	 			"01111110" 	when "01011111110",--6
				"00000000"	when "01011111111",--7
				--SPACE
				"00000000" 	when "00100000000",--0
				"00000000" 	when "00100000001",--1
				"00000000" 	when "00100000010",--2
				"00000000" 	when "00100000011",--3
				"00000000" 	when "00100000100",--4
				"00000000" 	when "00100000101",--5
	 			"00000000" 	when "00100000110",--6
				"00000000"	when "00100000111",--7
				--!
				"00011000" 	when "00100001000",--0
				"00011000" 	when "00100001001",--1
				"00011000" 	when "00100001010",--2
				"00011000" 	when "00100001011",--3
				"00000000" 	when "00100001100",--4
				"00000000" 	when "00100001101",--5
	 			"00011000" 	when "00100001110",--6
				"00000000"	when "00100001111",--7
				--"
				"01100110" 	when "00100010000",--0
				"01100110" 	when "00100010001",--1
				"01100110" 	when "00100010010",--2
				"00000000" 	when "00100010011",--3
				"00000000" 	when "00100010100",--4
				"00000000" 	when "00100010101",--5
	 			"00000000" 	when "00100010110",--6
				"00000000"	when "00100010111",--7
				--#
				"01100110" 	when "00100011000",--0
				"01100110" 	when "00100011001",--1
				"11111111" 	when "00100011010",--2
				"01100110" 	when "00100011011",--3
				"11111111" 	when "00100011100",--4
				"01100110" 	when "00100011101",--5
	 			"01100110" 	when "00100011110",--6
				"00000000"	when "00100011111",--7
				--$
				"00011000" 	when "00100100000",--0
				"00111110" 	when "00100100001",--1
				"01100000" 	when "00100100010",--2
				"00111100" 	when "00100100011",--3
				"00000110" 	when "00100100100",--4
				"01111100" 	when "00100100101",--5
	 			"00011000" 	when "00100100110",--6
				"00000000"	when "00100100111",--7
				--%
				"01100010" 	when "00100101000",--0
				"01100110" 	when "00100101001",--1
				"00001100" 	when "00100101010",--2
				"00011000" 	when "00100101011",--3
				"00110000" 	when "00100101100",--4
				"01100110" 	when "00100101101",--5
	 			"01000110" 	when "00100101110",--6
				"00000000"	when "00100101111",--7
				--&
				"00111100" 	when "00100110000",--0
				"01100110" 	when "00100110001",--1
				"00111100" 	when "00100110010",--2
				"00111000" 	when "00100110011",--3
				"01100111" 	when "00100110100",--4
				"01100110" 	when "00100110101",--5
	 			"00111111" 	when "00100110110",--6
				"00000000"	when "00100110111",--7
				--'
				"00000110" 	when "00100111000",--0
				"00001100" 	when "00100111001",--1
				"00011000" 	when "00100111010",--2
				"00000000" 	when "00100111011",--3
				"00000000" 	when "00100111100",--4
				"00000000" 	when "00100111101",--5
	 			"00000000" 	when "00100111110",--6
				"00000000"	when "00100111111",--7
				--(
				"00001100" 	when "00101000000",--0
				"00011000" 	when "00101000001",--1
				"00110000" 	when "00101000010",--2
				"00110000" 	when "00101000011",--3
				"00110000" 	when "00101000100",--4
				"00011000" 	when "00101000101",--5
	 			"00001100" 	when "00101000110",--6
				"00000000"	when "00101000111",--7
				--)
				"00110000" 	when "00101001000",--0
				"00011000" 	when "00101001001",--1
				"00001100" 	when "00101001010",--2
				"00001100" 	when "00101001011",--3
				"00001100" 	when "00101001100",--4
				"00011000" 	when "00101001101",--5
	 			"00110000" 	when "00101001110",--6
				"00000000"	when "00101001111",--7
				--*
				"00000000" 	when "00101010000",--0
				"01100110" 	when "00101010001",--1
				"00111100" 	when "00101010010",--2
				"11111111" 	when "00101010011",--3
				"00111100" 	when "00101010100",--4
				"01100110" 	when "00101010101",--5
	 			"00000000" 	when "00101010110",--6
				"00000000"	when "00101010111",--7
				--+
				"00000000" 	when "00101011000",--0
				"00011000" 	when "00101011001",--1
				"00011000" 	when "00101011010",--2
				"01111110" 	when "00101011011",--3
				"00011000" 	when "00101011100",--4
				"00011000" 	when "00101011101",--5
	 			"00000000" 	when "00101011110",--6
				"00000000"	when "00101011111",--7
				--,
				"00000000" 	when "00101100000",--0
				"00000000" 	when "00101100001",--1
				"00000000" 	when "00101100010",--2
				"00000000" 	when "00101100011",--3
				"00000000" 	when "00101100100",--4
				"00011000" 	when "00101100101",--5
	 			"00011000" 	when "00101100110",--6
				"00110000"	when "00101100111",--7
				---
				"00000000" 	when "00101101000",--0
				"00000000" 	when "00101101001",--1
				"00000000" 	when "00101101010",--2
				"01111110" 	when "00101101011",--3
				"00000000" 	when "00101101100",--4
				"00000000" 	when "00101101101",--5
	 			"00000000" 	when "00101101110",--6
				"00000000"	when "00101101111",--7
				--.
				"00000000" 	when "00101110000",--0
				"00000000" 	when "00101110001",--1
				"00000000" 	when "00101110010",--2
				"00000000" 	when "00101110011",--3
				"00000000" 	when "00101110100",--4
				"00000000" 	when "00101110101",--5
	 			"00011000" 	when "00101110110",--6
				"00000000"	when "00101110111",--7
				--/
				"00000000" 	when "00101111000",--0
				"00000011" 	when "00101111001",--1
				"00000110" 	when "00101111010",--2
				"00001100" 	when "00101111011",--3
				"00011000" 	when "00101111100",--4
				"00110000" 	when "00101111101",--5
	 			"01100000" 	when "00101111110",--6
				"00000000"	when "00101111111",--7
				--0
				"00111100" 	when "00110000000",--0
				"01100110" 	when "00110000001",--1
				"01101110" 	when "00110000010",--2
				"01110110" 	when "00110000011",--3
				"01100110" 	when "00110000100",--4
				"01100110" 	when "00110000101",--5
	 			"00111100" 	when "00110000110",--6
				"00000000"	when "00110000111",--7
				--1
				"00011000" 	when "00110001000",--0
				"00011000" 	when "00110001001",--1
				"00111000" 	when "00110001010",--2
				"00011000" 	when "00110001011",--3
				"00011000" 	when "00110001100",--4
				"00011000" 	when "00110001101",--5
	 			"01111110" 	when "00110001110",--6
				"00000000"	when "00110001111",--7
				--2
				"00111100" 	when "00110010000",--0
				"01100110" 	when "00110010001",--1
				"00000110" 	when "00110010010",--2
				"00001100" 	when "00110010011",--3
				"00110000" 	when "00110010100",--4
				"01100000" 	when "00110010101",--5
	 			"01111110" 	when "00110010110",--6
				"00000000"	when "00110010111",--7
				--3
				"00111100" 	when "00110011000",--0
				"01100110" 	when "00110011001",--1
				"00000110" 	when "00110011010",--2
				"00011100" 	when "00110011011",--3
				"00000110" 	when "00110011100",--4
				"01100110" 	when "00110011101",--5
	 			"00111100" 	when "00110011110",--6
				"00000000"	when "00110011111",--7
				--4
				"00000110" 	when "00110100000",--0
				"00001110" 	when "00110100001",--1
				"00011110" 	when "00110100010",--2
				"01100110" 	when "00110100011",--3
				"01111111" 	when "00110100100",--4
				"00000110" 	when "00110100101",--5
	 			"00000110" 	when "00110100110",--6
				"00000000"	when "00110100111",--7
				--5
				"01111110" 	when "00110101000",--0
				"01100000" 	when "00110101001",--1
				"01111100" 	when "00110101010",--2
				"00000110" 	when "00110101011",--3
				"00000110" 	when "00110101100",--4
				"01100110" 	when "00110101101",--5
	 			"00111100" 	when "00110101110",--6
				"00000000"	when "00110101111",--7
				--6
				"00111100" 	when "00110110000",--0
				"01100110" 	when "00110110001",--1
				"01100000" 	when "00110110010",--2
				"01111100" 	when "00110110011",--3
				"01100110" 	when "00110110100",--4
				"01100110" 	when "00110110101",--5
	 			"00111100" 	when "00110110110",--6
				"00000000"	when "00110110111",--7
				--7
				"01111110" 	when "00110111000",--0
				"01100110" 	when "00110111001",--1
				"00001100" 	when "00110111010",--2
				"00011000" 	when "00110111011",--3
				"00011000" 	when "00110111100",--4
				"00011000" 	when "00110111101",--5
	 			"00011000" 	when "00110111110",--6
				"00000000"	when "00110111111",--7
				--8
				"00111100" 	when "00111000000",--0
				"01100110" 	when "00111000001",--1
				"01100110" 	when "00111000010",--2
				"00111100" 	when "00111000011",--3
				"01100110" 	when "00111000100",--4
				"01100110" 	when "00111000101",--5
	 			"00111100" 	when "00111000110",--6
				"00000000"	when "00111000111",--7
				--9
				"00111100" 	when "00111001000",--0
				"01100110" 	when "00111001001",--1
				"01100110" 	when "00111001010",--2
				"00111110" 	when "00111001011",--3
				"00000110" 	when "00111001100",--4
				"01100110" 	when "00111001101",--5
	 			"00111100" 	when "00111001110",--6
				"00000000"	when "00111001111",--7
				--:
				"00000000" 	when "00111010000",--0
				"00000000" 	when "00111010001",--1
				"01100000" 	when "00111010010",--2
				"01100000" 	when "00111010011",--3
				"00000000" 	when "00111010100",--4
				"01100000" 	when "00111010101",--5
	 			"01100000" 	when "00111010110",--6
				"00000000"	when "00111010111",--7
				--;
				"00000000" 	when "00111011000",--0
				"00000000" 	when "00111011001",--1
				"01100000" 	when "00111011010",--2
				"01100000" 	when "00111011011",--3
				"00000000" 	when "00111011100",--4
				"01100000" 	when "00111011101",--5
	 			"01100000" 	when "00111011110",--6
				"11000000"	when "00111011111",--7
				--<
				"00000000" 	when "00111100000",--0
				"00000110" 	when "00111100001",--1
				"00011000" 	when "00111100010",--2
				"01100000" 	when "00111100011",--3
				"00011000" 	when "00111100100",--4
				"00000110" 	when "00111100101",--5
	 			"00000000" 	when "00111100110",--6
				"00000000"	when "00111100111",--7
				--=
				"00000000" 	when "00111101000",--0
				"00000000" 	when "00111101001",--1
				"01111110" 	when "00111101010",--2
				"00000000" 	when "00111101011",--3
				"01111110" 	when "00111101100",--4
				"00000000" 	when "00111101101",--5
	 			"00000000" 	when "00111101110",--6
				"00000000"	when "00111101111",--7
				-->
				"00000000" 	when "00111110000",--0
				"01100000" 	when "00111110001",--1
				"00011000" 	when "00111110010",--2
				"00000110" 	when "00111110011",--3
				"00011000" 	when "00111110100",--4
				"01100000" 	when "00111110101",--5
	 			"00000000" 	when "00111110110",--6
				"00000000"	when "00111110111",--7
				--?
				"00111100" 	when "00111111000",--0
				"11000110" 	when "00111111001",--1
				"00000110" 	when "00111111010",--2
				"00001100" 	when "00111111011",--3
				"00011000" 	when "00111111100",--4
				"00000000" 	when "00111111101",--5
	 			"00011000" 	when "00111111110",--6
				"00000000"	when "00111111111",--7
				--`
				"01100000" 	when "01100000000",
				"00110000" 	when "01100000001",
				"00011000" 	when "01100000010",
				"00000000" 	when "01100000011",
				"00000000" 	when "01100000100",
				"00000000" 	when "01100000101",
	 			"00000000" 	when "01100000110",
				"00000000" 	when "01100000111",
				--a
				"00000000"	when "01100001000",
				"00000000"	when "01100001001",
				"00111100"	when "01100001010",
				"00000110"	when "01100001011",
				"00111110"	when "01100001100",
				"01100110"	when "01100001101",
				"00111110"	when "01100001110",
				"00000000"	when "01100001111",
				--b
				"01100000" 	when "01100010000",
				"01100000" 	when "01100010001",
				"01111100" 	when "01100010010",
				"01100110" 	when "01100010011",
				"01100110" 	when "01100010100",
				"01100110" 	when "01100010101",
	 			"01111100" 	when "01100010110",
				"00000000"	when "01100010111",				

				--c
				"00000000" 	when "01100011000",
				"00000000" 	when "01100011001",
				"00111100" 	when "01100011010",
				"01100110" 	when "01100011011",
				"01100000" 	when "01100011100",
				"01100110" 	when "01100011101",
	 			"00111100" 	when "01100011110",
				"00000000"	when "01100011111",
				--d
				"00000110" 	when "01100100000",
				"00000110" 	when "01100100001",
				"00111110" 	when "01100100010",
				"01100110" 	when "01100100011",
				"01100110" 	when "01100100100",
				"01100110" 	when "01100100101",
	 			"00111110" 	when "01100100110",
				"00000000"	when "01100100111",				

				--e
				"00000000" 	when "01100101000",
				"00000000" 	when "01100101001",
				"00111100" 	when "01100101010",
				"01100110" 	when "01100101011",
				"01111110" 	when "01100101100",
				"01100000" 	when "01100101101",
	 			"00111110" 	when "01100101110",
				"00000000"	when "01100101111",
				--f
				"00011100" 	when "01100110000",--0
				"00110000" 	when "01100110001",--1
				"00110000" 	when "01100110010",--2
				"01111100" 	when "01100110011",--3
				"00110000" 	when "01100110100",--4
				"00110000" 	when "01100110101",--5
	 			"00110000" 	when "01100110110",--6
				"00000000"	when "01100110111",--7
				--g
				"00000000" 	when "01100111000",--0
				"00000000" 	when "01100111001",--1
				"00111110" 	when "01100111010",--2
				"01100110" 	when "01100111011",--3
				"01100110" 	when "01100111100",--4
				"00111110" 	when "01100111101",--5
	 			"00000110" 	when "01100111110",--6
				"01111100"	when "01100111111",--7
				--h
				"01100000" 	when "01101000000",--0
				"01100000" 	when "01101000001",--1
				"01111100" 	when "01101000010",--2
				"01100110" 	when "01101000011",--3
				"01100110" 	when "01101000100",--4
				"01100110" 	when "01101000101",--5
	 			"01100110" 	when "01101000110",--6
				"00000000"	when "01101000111",--7
				--i
				"00011000" 	when "01101001000",--0
				"00000000" 	when "01101001001",--1
				"00011000" 	when "01101001010",--2
				"00011000" 	when "01101001011",--3
				"00011000" 	when "01101001100",--4
				"00011000" 	when "01101001101",--5
	 			"00011000" 	when "01101001110",--6
				"00000000"	when "01101001111",--7
				--j
				"00001100" 	when "01101010000",--0
				"00000000" 	when "01101010001",--1
				"00001100" 	when "01101010010",--2
				"00001100" 	when "01101010011",--3
				"00001100" 	when "01101010100",--4
				"00001100" 	when "01101010101",--5
	 			"01101100" 	when "01101010110",--6
				"00111000"	when "01101010111",--7
				--k
				"01100000" 	when "01101011000",--0
				"01100000" 	when "01101011001",--1
				"01100110" 	when "01101011010",--2
				"01101100" 	when "01101011011",--3
				"01111000" 	when "01101011100",--4
				"01101100" 	when "01101011101",--5
	 			"01100110" 	when "01101011110",--6
				"00000000"	when "01101011111",--7
				--l
				"00111000" 	when "01101100000",--0
				"00011000" 	when "01101100001",--1
				"00011000" 	when "01101100010",--2
				"00011000" 	when "01101100011",--3
				"00011000" 	when "01101100100",--4
				"00011000" 	when "01101100101",--5
	 			"00111100" 	when "01101100110",--6
				"00000000"	when "01101100111",--7
				--m
				"00000000" 	when "01101101000",--0
				"00000000" 	when "01101101001",--1
				"11110110" 	when "01101101010",--2
				"11011011" 	when "01101101011",--3
				"11011011" 	when "01101101100",--4
				"11011011" 	when "01101101101",--5
	 			"11011011" 	when "01101101110",--6
				"00000000"	when "01101101111",--7
				--n
				"00000000" 	when "01101110000",--0
				"00000000" 	when "01101110001",--1
				"01111100" 	when "01101110010",--2
				"01100110" 	when "01101110011",--3
				"01100110" 	when "01101110100",--4
				"01100110" 	when "01101110101",--5
	 			"01100110" 	when "01101110110",--6
				"00000000"	when "01101110111",--7
				--o
				"00000000" 	when "01101111000",--0
				"00000000" 	when "01101111001",--1
				"00111100" 	when "01101111010",--2
				"01100110" 	when "01101111011",--3
				"01100110" 	when "01101111100",--4
				"01100110" 	when "01101111101",--5
	 			"00111100" 	when "01101111110",--6
				"00000000"	when "01101111111",--7
				--p
				"00000000" 	when "01110000000",--0
				"00000000" 	when "01110000001",--1
				"01111100" 	when "01110000010",--2
				"01100110" 	when "01110000011",--3
				"01100110" 	when "01110000100",--4
				"01111100" 	when "01110000101",--5
	 			"01100000" 	when "01110000110",--6
				"01100000"	when "01110000111",--7
				--q
				"00000000" 	when "01110001000",--0
				"00000000" 	when "01110001001",--1
				"00111110" 	when "01110001010",--2
				"01100110" 	when "01110001011",--3
				"01100110" 	when "01110001100",--4
				"00111110" 	when "01110001101",--5
	 			"00000110" 	when "01110001110",--6
				"00000110"	when "01110001111",--7
				--r
				"00000000" 	when "01110010000",--0
				"00000000" 	when "01110010001",--1
				"01101100" 	when "01110010010",--2
				"01111000" 	when "01110010011",--3
				"01100000" 	when "01110010100",--4
				"01100000" 	when "01110010101",--5
	 			"01100000" 	when "01110010110",--6
				"00000000"	when "01110010111",--7
				--s
				"00000000" 	when "01110011000",--0
				"00000000" 	when "01110011001",--1
				"00111110" 	when "01110011010",--2
				"01100000" 	when "01110011011",--3
				"00111100" 	when "01110011100",--4
				"00000110" 	when "01110011101",--5
	 			"01111100" 	when "01110011110",--6
				"00000000"	when "01110011111",--7
				--t
				"00000000" 	when "01110100000",--0
				"00110000" 	when "01110100001",--1
				"01111100" 	when "01110100010",--2
				"00110000" 	when "01110100011",--3
				"00110000" 	when "01110100100",--4
				"00110000" 	when "01110100101",--5
	 			"00011100" 	when "01110100110",--6
				"00000000"	when "01110100111",--7
				--u
				"00000000" 	when "01110101000",--0
				"00000000" 	when "01110101001",--1
				"01100110" 	when "01110101010",--2
				"01100110" 	when "01110101011",--3
				"01100110" 	when "01110101100",--4
				"01100110" 	when "01110101101",--5
	 			"00111110" 	when "01110101110",--6
				"00000000"	when "01110101111",--7
				--v
				"00000000" 	when "01110110000",--0
				"00000000" 	when "01110110001",--1
				"01100110" 	when "01110110010",--2
				"01100110" 	when "01110110011",--3
				"01100110" 	when "01110110100",--4
				"00111100" 	when "01110110101",--5
	 			"00011000" 	when "01110110110",--6
				"00000000"	when "01110110111",--7
				--w
				"00000000" 	when "01110111000",--0
				"00000000" 	when "01110111001",--1
				"11000011" 	when "01110111010",--2
				"11000011" 	when "01110111011",--3
				"11011011" 	when "01110111100",--4
				"11011011" 	when "01110111101",--5
	 			"01100110" 	when "01110111110",--6
				"00000000"	when "01110111111",--7
				--x
				"00000000" 	when "01111000000",--0
				"00000000" 	when "01111000001",--1
				"01100110" 	when "01111000010",--2
				"00011000" 	when "01111000011",--3
				"00011000" 	when "01111000100",--4
				"00011000" 	when "01111000101",--5
	 			"01100110" 	when "01111000110",--6
				"00000000"	when "01111000111",--7
				--y
				"00000000" 	when "01111001000",--0
				"00000000" 	when "01111001001",--1
				"01100110" 	when "01111001010",--2
				"01100110" 	when "01111001011",--3
				"01100110" 	when "01111001100",--4
				"00111110" 	when "01111001101",--5
	 			"00000110" 	when "01111001110",--6
				"00111100"	when "01111001111",--7
				--z
				"00000000" 	when "01111010000",--0
				"00000000" 	when "01111010001",--1
				"01111110" 	when "01111010010",--2
				"00001100" 	when "01111010011",--3
				"00011000" 	when "01111010100",--4
				"00110000" 	when "01111010101",--5
	 			"01111110" 	when "01111010110",--6
				"00000000"	when "01111010111",--7
				--{
				"00011000" 	when "01111011000",--0
				"00110000" 	when "01111011001",--1
				"00110000" 	when "01111011010",--2
				"01110000" 	when "01111011011",--3
				"00110000" 	when "01111011100",--4
				"00110000" 	when "01111011101",--5
	 			"00011000" 	when "01111011110",--6
				"00000000"	when "01111011111",--7
				--|
				"00011000" 	when "01111100000",--0
				"00011000" 	when "01111100001",--1
				"00011000" 	when "01111100010",--2
				"00011000" 	when "01111100011",--3
				"00011000" 	when "01111100100",--4
				"00011000" 	when "01111100101",--5
	 			"00011000" 	when "01111100110",--6
				"00000000"	when "01111100111",--7
				--}
				"00011000" 	when "01111101000",--0
				"00001100" 	when "01111101001",--1
				"00001100" 	when "01111101010",--2
				"00001110" 	when "01111101011",--3
				"00001100" 	when "01111101100",--4
				"00001100" 	when "01111101101",--5
	 			"00011000" 	when "01111101110",--6
				"00000000"	when "01111101111",--7
				--~
				"00000000" 	when "01111110000",--0
				"00000000" 	when "01111110001",--1
				"01110000" 	when "01111110010",--2
				"11011011" 	when "01111110011",--3
				"00001110" 	when "01111110100",--4
				"00000000" 	when "01111110101",--5
	 			"00000000" 	when "01111110110",--6
				"00000000"	when "01111110111",--7
				-- 
				"00000000"	when others;
				
				


rom_address <= character_address & font_row;

rom_mux_output <= rom_data ( (CONV_INTEGER(NOT font_col(2 DOWNTO 0))));

END a;